module layer0_N116 ( input [6:0] M0, output [1:0] M1 );

	(*rom_style = "distributed" *) reg [1:0] M1r;
	assign M1 = M1r;
	always @ (M0) begin
		case (M0)
			7'b0000000: M1r = 2'b00;
			7'b1000000: M1r = 2'b00;
			7'b0100000: M1r = 2'b00;
			7'b1100000: M1r = 2'b00;
			7'b0010000: M1r = 2'b00;
			7'b1010000: M1r = 2'b00;
			7'b0110000: M1r = 2'b00;
			7'b1110000: M1r = 2'b00;
			7'b0001000: M1r = 2'b00;
			7'b1001000: M1r = 2'b01;
			7'b0101000: M1r = 2'b00;
			7'b1101000: M1r = 2'b00;
			7'b0011000: M1r = 2'b00;
			7'b1011000: M1r = 2'b01;
			7'b0111000: M1r = 2'b00;
			7'b1111000: M1r = 2'b00;
			7'b0000100: M1r = 2'b00;
			7'b1000100: M1r = 2'b01;
			7'b0100100: M1r = 2'b00;
			7'b1100100: M1r = 2'b00;
			7'b0010100: M1r = 2'b00;
			7'b1010100: M1r = 2'b01;
			7'b0110100: M1r = 2'b00;
			7'b1110100: M1r = 2'b00;
			7'b0001100: M1r = 2'b10;
			7'b1001100: M1r = 2'b10;
			7'b0101100: M1r = 2'b01;
			7'b1101100: M1r = 2'b10;
			7'b0011100: M1r = 2'b10;
			7'b1011100: M1r = 2'b10;
			7'b0111100: M1r = 2'b01;
			7'b1111100: M1r = 2'b01;
			7'b0000010: M1r = 2'b00;
			7'b1000010: M1r = 2'b00;
			7'b0100010: M1r = 2'b00;
			7'b1100010: M1r = 2'b00;
			7'b0010010: M1r = 2'b00;
			7'b1010010: M1r = 2'b00;
			7'b0110010: M1r = 2'b00;
			7'b1110010: M1r = 2'b00;
			7'b0001010: M1r = 2'b01;
			7'b1001010: M1r = 2'b10;
			7'b0101010: M1r = 2'b01;
			7'b1101010: M1r = 2'b01;
			7'b0011010: M1r = 2'b01;
			7'b1011010: M1r = 2'b10;
			7'b0111010: M1r = 2'b00;
			7'b1111010: M1r = 2'b01;
			7'b0000110: M1r = 2'b01;
			7'b1000110: M1r = 2'b10;
			7'b0100110: M1r = 2'b00;
			7'b1100110: M1r = 2'b01;
			7'b0010110: M1r = 2'b01;
			7'b1010110: M1r = 2'b01;
			7'b0110110: M1r = 2'b00;
			7'b1110110: M1r = 2'b01;
			7'b0001110: M1r = 2'b11;
			7'b1001110: M1r = 2'b11;
			7'b0101110: M1r = 2'b10;
			7'b1101110: M1r = 2'b11;
			7'b0011110: M1r = 2'b10;
			7'b1011110: M1r = 2'b11;
			7'b0111110: M1r = 2'b10;
			7'b1111110: M1r = 2'b10;
			7'b0000001: M1r = 2'b00;
			7'b1000001: M1r = 2'b00;
			7'b0100001: M1r = 2'b00;
			7'b1100001: M1r = 2'b00;
			7'b0010001: M1r = 2'b00;
			7'b1010001: M1r = 2'b00;
			7'b0110001: M1r = 2'b00;
			7'b1110001: M1r = 2'b00;
			7'b0001001: M1r = 2'b00;
			7'b1001001: M1r = 2'b00;
			7'b0101001: M1r = 2'b00;
			7'b1101001: M1r = 2'b00;
			7'b0011001: M1r = 2'b00;
			7'b1011001: M1r = 2'b00;
			7'b0111001: M1r = 2'b00;
			7'b1111001: M1r = 2'b00;
			7'b0000101: M1r = 2'b00;
			7'b1000101: M1r = 2'b00;
			7'b0100101: M1r = 2'b00;
			7'b1100101: M1r = 2'b00;
			7'b0010101: M1r = 2'b00;
			7'b1010101: M1r = 2'b00;
			7'b0110101: M1r = 2'b00;
			7'b1110101: M1r = 2'b00;
			7'b0001101: M1r = 2'b00;
			7'b1001101: M1r = 2'b01;
			7'b0101101: M1r = 2'b00;
			7'b1101101: M1r = 2'b00;
			7'b0011101: M1r = 2'b00;
			7'b1011101: M1r = 2'b01;
			7'b0111101: M1r = 2'b00;
			7'b1111101: M1r = 2'b00;
			7'b0000011: M1r = 2'b00;
			7'b1000011: M1r = 2'b00;
			7'b0100011: M1r = 2'b00;
			7'b1100011: M1r = 2'b00;
			7'b0010011: M1r = 2'b00;
			7'b1010011: M1r = 2'b00;
			7'b0110011: M1r = 2'b00;
			7'b1110011: M1r = 2'b00;
			7'b0001011: M1r = 2'b00;
			7'b1001011: M1r = 2'b01;
			7'b0101011: M1r = 2'b00;
			7'b1101011: M1r = 2'b00;
			7'b0011011: M1r = 2'b00;
			7'b1011011: M1r = 2'b00;
			7'b0111011: M1r = 2'b00;
			7'b1111011: M1r = 2'b00;
			7'b0000111: M1r = 2'b00;
			7'b1000111: M1r = 2'b00;
			7'b0100111: M1r = 2'b00;
			7'b1100111: M1r = 2'b00;
			7'b0010111: M1r = 2'b00;
			7'b1010111: M1r = 2'b00;
			7'b0110111: M1r = 2'b00;
			7'b1110111: M1r = 2'b00;
			7'b0001111: M1r = 2'b01;
			7'b1001111: M1r = 2'b10;
			7'b0101111: M1r = 2'b00;
			7'b1101111: M1r = 2'b01;
			7'b0011111: M1r = 2'b01;
			7'b1011111: M1r = 2'b10;
			7'b0111111: M1r = 2'b00;
			7'b1111111: M1r = 2'b01;

		endcase
	end
endmodule

module layer0 (input [47:0] M0, output [144:0] M1);

wire [5:0] layer0_N0_wire = {M0[47], M0[45], M0[35], M0[30], M0[15], M0[7]};
layer0_N0 layer0_N0_inst (.M0(layer0_N0_wire), .M1(M1[0:0]));

wire [5:0] layer0_N1_wire = {M0[40], M0[34], M0[19], M0[16], M0[9], M0[7]};
layer0_N1 layer0_N1_inst (.M0(layer0_N1_wire), .M1(M1[1:1]));

wire [5:0] layer0_N2_wire = {M0[31], M0[21], M0[15], M0[14], M0[12], M0[9]};
layer0_N2 layer0_N2_inst (.M0(layer0_N2_wire), .M1(M1[2:2]));

wire [5:0] layer0_N3_wire = {M0[36], M0[34], M0[24], M0[13], M0[12], M0[1]};
layer0_N3 layer0_N3_inst (.M0(layer0_N3_wire), .M1(M1[3:3]));

wire [5:0] layer0_N4_wire = {M0[47], M0[43], M0[35], M0[27], M0[24], M0[8]};
layer0_N4 layer0_N4_inst (.M0(layer0_N4_wire), .M1(M1[4:4]));

wire [5:0] layer0_N5_wire = {M0[45], M0[38], M0[28], M0[27], M0[24], M0[0]};
layer0_N5 layer0_N5_inst (.M0(layer0_N5_wire), .M1(M1[5:5]));

wire [5:0] layer0_N6_wire = {M0[45], M0[40], M0[34], M0[21], M0[18], M0[13]};
layer0_N6 layer0_N6_inst (.M0(layer0_N6_wire), .M1(M1[6:6]));

wire [5:0] layer0_N7_wire = {M0[47], M0[40], M0[30], M0[23], M0[14], M0[10]};
layer0_N7 layer0_N7_inst (.M0(layer0_N7_wire), .M1(M1[7:7]));

wire [5:0] layer0_N8_wire = {M0[38], M0[37], M0[18], M0[10], M0[4], M0[1]};
layer0_N8 layer0_N8_inst (.M0(layer0_N8_wire), .M1(M1[8:8]));

wire [5:0] layer0_N9_wire = {M0[43], M0[28], M0[11], M0[6], M0[2], M0[0]};
layer0_N9 layer0_N9_inst (.M0(layer0_N9_wire), .M1(M1[9:9]));

wire [5:0] layer0_N10_wire = {M0[45], M0[39], M0[38], M0[29], M0[16], M0[3]};
layer0_N10 layer0_N10_inst (.M0(layer0_N10_wire), .M1(M1[10:10]));

wire [5:0] layer0_N11_wire = {M0[28], M0[23], M0[20], M0[14], M0[9], M0[0]};
layer0_N11 layer0_N11_inst (.M0(layer0_N11_wire), .M1(M1[11:11]));

wire [5:0] layer0_N12_wire = {M0[47], M0[46], M0[30], M0[26], M0[24], M0[2]};
layer0_N12 layer0_N12_inst (.M0(layer0_N12_wire), .M1(M1[12:12]));

wire [5:0] layer0_N13_wire = {M0[40], M0[35], M0[34], M0[32], M0[29], M0[10]};
layer0_N13 layer0_N13_inst (.M0(layer0_N13_wire), .M1(M1[13:13]));

wire [5:0] layer0_N14_wire = {M0[44], M0[42], M0[31], M0[21], M0[12], M0[1]};
layer0_N14 layer0_N14_inst (.M0(layer0_N14_wire), .M1(M1[14:14]));

wire [5:0] layer0_N15_wire = {M0[45], M0[37], M0[31], M0[12], M0[7], M0[3]};
layer0_N15 layer0_N15_inst (.M0(layer0_N15_wire), .M1(M1[15:15]));

wire [5:0] layer0_N16_wire = {M0[37], M0[33], M0[27], M0[21], M0[15], M0[11]};
layer0_N16 layer0_N16_inst (.M0(layer0_N16_wire), .M1(M1[16:16]));

wire [5:0] layer0_N17_wire = {M0[38], M0[30], M0[23], M0[17], M0[14], M0[0]};
layer0_N17 layer0_N17_inst (.M0(layer0_N17_wire), .M1(M1[17:17]));

wire [5:0] layer0_N18_wire = {M0[24], M0[22], M0[19], M0[15], M0[9], M0[4]};
layer0_N18 layer0_N18_inst (.M0(layer0_N18_wire), .M1(M1[18:18]));

wire [5:0] layer0_N19_wire = {M0[36], M0[31], M0[26], M0[20], M0[18], M0[10]};
layer0_N19 layer0_N19_inst (.M0(layer0_N19_wire), .M1(M1[19:19]));

wire [5:0] layer0_N20_wire = {M0[40], M0[38], M0[20], M0[11], M0[4], M0[1]};
layer0_N20 layer0_N20_inst (.M0(layer0_N20_wire), .M1(M1[20:20]));

wire [5:0] layer0_N21_wire = {M0[45], M0[34], M0[24], M0[16], M0[5], M0[0]};
layer0_N21 layer0_N21_inst (.M0(layer0_N21_wire), .M1(M1[21:21]));

wire [5:0] layer0_N22_wire = {M0[44], M0[38], M0[29], M0[26], M0[18], M0[9]};
layer0_N22 layer0_N22_inst (.M0(layer0_N22_wire), .M1(M1[22:22]));

wire [5:0] layer0_N23_wire = {M0[47], M0[41], M0[37], M0[26], M0[6], M0[2]};
layer0_N23 layer0_N23_inst (.M0(layer0_N23_wire), .M1(M1[23:23]));

wire [5:0] layer0_N24_wire = {M0[38], M0[37], M0[35], M0[33], M0[15], M0[11]};
layer0_N24 layer0_N24_inst (.M0(layer0_N24_wire), .M1(M1[24:24]));

wire [5:0] layer0_N25_wire = {M0[40], M0[35], M0[32], M0[30], M0[9], M0[1]};
layer0_N25 layer0_N25_inst (.M0(layer0_N25_wire), .M1(M1[25:25]));

wire [5:0] layer0_N26_wire = {M0[47], M0[30], M0[25], M0[9], M0[7], M0[1]};
layer0_N26 layer0_N26_inst (.M0(layer0_N26_wire), .M1(M1[26:26]));

wire [5:0] layer0_N27_wire = {M0[46], M0[27], M0[25], M0[16], M0[8], M0[4]};
layer0_N27 layer0_N27_inst (.M0(layer0_N27_wire), .M1(M1[27:27]));

wire [5:0] layer0_N28_wire = {M0[29], M0[28], M0[25], M0[24], M0[14], M0[12]};
layer0_N28 layer0_N28_inst (.M0(layer0_N28_wire), .M1(M1[28:28]));

wire [5:0] layer0_N29_wire = {M0[26], M0[25], M0[22], M0[14], M0[11], M0[8]};
layer0_N29 layer0_N29_inst (.M0(layer0_N29_wire), .M1(M1[29:29]));

wire [5:0] layer0_N30_wire = {M0[45], M0[29], M0[27], M0[12], M0[11], M0[8]};
layer0_N30 layer0_N30_inst (.M0(layer0_N30_wire), .M1(M1[30:30]));

wire [5:0] layer0_N31_wire = {M0[45], M0[33], M0[30], M0[28], M0[19], M0[5]};
layer0_N31 layer0_N31_inst (.M0(layer0_N31_wire), .M1(M1[31:31]));

wire [5:0] layer0_N32_wire = {M0[43], M0[40], M0[32], M0[11], M0[7], M0[3]};
layer0_N32 layer0_N32_inst (.M0(layer0_N32_wire), .M1(M1[32:32]));

wire [5:0] layer0_N33_wire = {M0[40], M0[19], M0[15], M0[8], M0[7], M0[3]};
layer0_N33 layer0_N33_inst (.M0(layer0_N33_wire), .M1(M1[33:33]));

wire [5:0] layer0_N34_wire = {M0[40], M0[33], M0[31], M0[21], M0[20], M0[8]};
layer0_N34 layer0_N34_inst (.M0(layer0_N34_wire), .M1(M1[34:34]));

wire [5:0] layer0_N35_wire = {M0[43], M0[34], M0[23], M0[18], M0[17], M0[15]};
layer0_N35 layer0_N35_inst (.M0(layer0_N35_wire), .M1(M1[35:35]));

wire [5:0] layer0_N36_wire = {M0[40], M0[39], M0[37], M0[36], M0[15], M0[11]};
layer0_N36 layer0_N36_inst (.M0(layer0_N36_wire), .M1(M1[36:36]));

wire [5:0] layer0_N37_wire = {M0[47], M0[46], M0[43], M0[42], M0[32], M0[6]};
layer0_N37 layer0_N37_inst (.M0(layer0_N37_wire), .M1(M1[37:37]));

wire [5:0] layer0_N38_wire = {M0[45], M0[34], M0[22], M0[21], M0[16], M0[10]};
layer0_N38 layer0_N38_inst (.M0(layer0_N38_wire), .M1(M1[38:38]));

wire [5:0] layer0_N39_wire = {M0[38], M0[33], M0[18], M0[10], M0[9], M0[6]};
layer0_N39 layer0_N39_inst (.M0(layer0_N39_wire), .M1(M1[39:39]));

wire [5:0] layer0_N40_wire = {M0[41], M0[29], M0[20], M0[19], M0[11], M0[7]};
layer0_N40 layer0_N40_inst (.M0(layer0_N40_wire), .M1(M1[40:40]));

wire [5:0] layer0_N41_wire = {M0[37], M0[34], M0[17], M0[13], M0[12], M0[0]};
layer0_N41 layer0_N41_inst (.M0(layer0_N41_wire), .M1(M1[41:41]));

wire [5:0] layer0_N42_wire = {M0[47], M0[39], M0[38], M0[14], M0[8], M0[4]};
layer0_N42 layer0_N42_inst (.M0(layer0_N42_wire), .M1(M1[42:42]));

wire [5:0] layer0_N43_wire = {M0[43], M0[37], M0[19], M0[8], M0[5], M0[3]};
layer0_N43 layer0_N43_inst (.M0(layer0_N43_wire), .M1(M1[43:43]));

wire [5:0] layer0_N44_wire = {M0[40], M0[34], M0[31], M0[30], M0[28], M0[5]};
layer0_N44 layer0_N44_inst (.M0(layer0_N44_wire), .M1(M1[44:44]));

wire [5:0] layer0_N45_wire = {M0[36], M0[33], M0[31], M0[13], M0[3], M0[0]};
layer0_N45 layer0_N45_inst (.M0(layer0_N45_wire), .M1(M1[45:45]));

wire [5:0] layer0_N46_wire = {M0[42], M0[29], M0[20], M0[18], M0[14], M0[7]};
layer0_N46 layer0_N46_inst (.M0(layer0_N46_wire), .M1(M1[46:46]));

wire [5:0] layer0_N47_wire = {M0[42], M0[38], M0[29], M0[28], M0[21], M0[12]};
layer0_N47 layer0_N47_inst (.M0(layer0_N47_wire), .M1(M1[47:47]));

wire [5:0] layer0_N48_wire = {M0[45], M0[36], M0[31], M0[27], M0[2], M0[1]};
layer0_N48 layer0_N48_inst (.M0(layer0_N48_wire), .M1(M1[48:48]));

wire [5:0] layer0_N49_wire = {M0[42], M0[37], M0[36], M0[29], M0[23], M0[6]};
layer0_N49 layer0_N49_inst (.M0(layer0_N49_wire), .M1(M1[49:49]));

wire [5:0] layer0_N50_wire = {M0[44], M0[37], M0[22], M0[4], M0[3], M0[1]};
layer0_N50 layer0_N50_inst (.M0(layer0_N50_wire), .M1(M1[50:50]));

wire [5:0] layer0_N51_wire = {M0[42], M0[39], M0[36], M0[29], M0[21], M0[10]};
layer0_N51 layer0_N51_inst (.M0(layer0_N51_wire), .M1(M1[51:51]));

wire [5:0] layer0_N52_wire = {M0[45], M0[44], M0[18], M0[13], M0[4], M0[3]};
layer0_N52 layer0_N52_inst (.M0(layer0_N52_wire), .M1(M1[52:52]));

wire [5:0] layer0_N53_wire = {M0[33], M0[29], M0[27], M0[18], M0[10], M0[8]};
layer0_N53 layer0_N53_inst (.M0(layer0_N53_wire), .M1(M1[53:53]));

wire [5:0] layer0_N54_wire = {M0[47], M0[37], M0[36], M0[32], M0[23], M0[14]};
layer0_N54 layer0_N54_inst (.M0(layer0_N54_wire), .M1(M1[54:54]));

wire [5:0] layer0_N55_wire = {M0[34], M0[32], M0[26], M0[18], M0[14], M0[5]};
layer0_N55 layer0_N55_inst (.M0(layer0_N55_wire), .M1(M1[55:55]));

wire [5:0] layer0_N56_wire = {M0[38], M0[29], M0[23], M0[11], M0[10], M0[5]};
layer0_N56 layer0_N56_inst (.M0(layer0_N56_wire), .M1(M1[56:56]));

wire [5:0] layer0_N57_wire = {M0[47], M0[41], M0[38], M0[28], M0[25], M0[15]};
layer0_N57 layer0_N57_inst (.M0(layer0_N57_wire), .M1(M1[57:57]));

wire [5:0] layer0_N58_wire = {M0[44], M0[43], M0[39], M0[28], M0[13], M0[4]};
layer0_N58 layer0_N58_inst (.M0(layer0_N58_wire), .M1(M1[58:58]));

wire [5:0] layer0_N59_wire = {M0[36], M0[32], M0[24], M0[8], M0[7], M0[0]};
layer0_N59 layer0_N59_inst (.M0(layer0_N59_wire), .M1(M1[59:59]));

wire [5:0] layer0_N60_wire = {M0[25], M0[24], M0[22], M0[15], M0[10], M0[6]};
layer0_N60 layer0_N60_inst (.M0(layer0_N60_wire), .M1(M1[60:60]));

wire [5:0] layer0_N61_wire = {M0[41], M0[31], M0[27], M0[15], M0[7], M0[2]};
layer0_N61 layer0_N61_inst (.M0(layer0_N61_wire), .M1(M1[61:61]));

wire [5:0] layer0_N62_wire = {M0[40], M0[37], M0[31], M0[24], M0[17], M0[13]};
layer0_N62 layer0_N62_inst (.M0(layer0_N62_wire), .M1(M1[62:62]));

wire [5:0] layer0_N63_wire = {M0[47], M0[42], M0[41], M0[37], M0[34], M0[33]};
layer0_N63 layer0_N63_inst (.M0(layer0_N63_wire), .M1(M1[63:63]));

wire [5:0] layer0_N64_wire = {M0[47], M0[46], M0[44], M0[30], M0[26], M0[12]};
layer0_N64 layer0_N64_inst (.M0(layer0_N64_wire), .M1(M1[64:64]));

wire [5:0] layer0_N65_wire = {M0[44], M0[37], M0[36], M0[29], M0[24], M0[12]};
layer0_N65 layer0_N65_inst (.M0(layer0_N65_wire), .M1(M1[65:65]));

wire [5:0] layer0_N66_wire = {M0[27], M0[26], M0[22], M0[21], M0[15], M0[13]};
layer0_N66 layer0_N66_inst (.M0(layer0_N66_wire), .M1(M1[66:66]));

wire [5:0] layer0_N67_wire = {M0[45], M0[43], M0[33], M0[22], M0[6], M0[0]};
layer0_N67 layer0_N67_inst (.M0(layer0_N67_wire), .M1(M1[67:67]));

wire [5:0] layer0_N68_wire = {M0[32], M0[30], M0[22], M0[18], M0[10], M0[0]};
layer0_N68 layer0_N68_inst (.M0(layer0_N68_wire), .M1(M1[68:68]));

wire [5:0] layer0_N69_wire = {M0[36], M0[30], M0[29], M0[24], M0[12], M0[8]};
layer0_N69 layer0_N69_inst (.M0(layer0_N69_wire), .M1(M1[69:69]));

wire [5:0] layer0_N70_wire = {M0[44], M0[35], M0[19], M0[17], M0[10], M0[1]};
layer0_N70 layer0_N70_inst (.M0(layer0_N70_wire), .M1(M1[70:70]));

wire [5:0] layer0_N71_wire = {M0[47], M0[41], M0[28], M0[19], M0[18], M0[2]};
layer0_N71 layer0_N71_inst (.M0(layer0_N71_wire), .M1(M1[71:71]));

wire [5:0] layer0_N72_wire = {M0[46], M0[43], M0[37], M0[24], M0[23], M0[6]};
layer0_N72 layer0_N72_inst (.M0(layer0_N72_wire), .M1(M1[72:72]));

wire [5:0] layer0_N73_wire = {M0[41], M0[37], M0[15], M0[10], M0[8], M0[3]};
layer0_N73 layer0_N73_inst (.M0(layer0_N73_wire), .M1(M1[73:73]));

wire [5:0] layer0_N74_wire = {M0[35], M0[32], M0[31], M0[28], M0[9], M0[5]};
layer0_N74 layer0_N74_inst (.M0(layer0_N74_wire), .M1(M1[74:74]));

wire [5:0] layer0_N75_wire = {M0[44], M0[41], M0[35], M0[22], M0[21], M0[17]};
layer0_N75 layer0_N75_inst (.M0(layer0_N75_wire), .M1(M1[75:75]));

wire [5:0] layer0_N76_wire = {M0[44], M0[43], M0[32], M0[18], M0[7], M0[2]};
layer0_N76 layer0_N76_inst (.M0(layer0_N76_wire), .M1(M1[76:76]));

wire [5:0] layer0_N77_wire = {M0[37], M0[22], M0[11], M0[10], M0[7], M0[6]};
layer0_N77 layer0_N77_inst (.M0(layer0_N77_wire), .M1(M1[77:77]));

wire [5:0] layer0_N78_wire = {M0[37], M0[35], M0[34], M0[27], M0[19], M0[7]};
layer0_N78 layer0_N78_inst (.M0(layer0_N78_wire), .M1(M1[78:78]));

wire [5:0] layer0_N79_wire = {M0[32], M0[23], M0[15], M0[14], M0[6], M0[5]};
layer0_N79 layer0_N79_inst (.M0(layer0_N79_wire), .M1(M1[79:79]));

wire [5:0] layer0_N80_wire = {M0[45], M0[36], M0[33], M0[24], M0[12], M0[0]};
layer0_N80 layer0_N80_inst (.M0(layer0_N80_wire), .M1(M1[80:80]));

wire [5:0] layer0_N81_wire = {M0[46], M0[25], M0[18], M0[8], M0[5], M0[4]};
layer0_N81 layer0_N81_inst (.M0(layer0_N81_wire), .M1(M1[81:81]));

wire [5:0] layer0_N82_wire = {M0[42], M0[29], M0[28], M0[24], M0[17], M0[3]};
layer0_N82 layer0_N82_inst (.M0(layer0_N82_wire), .M1(M1[82:82]));

wire [5:0] layer0_N83_wire = {M0[44], M0[33], M0[30], M0[27], M0[15], M0[5]};
layer0_N83 layer0_N83_inst (.M0(layer0_N83_wire), .M1(M1[83:83]));

wire [5:0] layer0_N84_wire = {M0[47], M0[44], M0[40], M0[37], M0[6], M0[3]};
layer0_N84 layer0_N84_inst (.M0(layer0_N84_wire), .M1(M1[84:84]));

wire [5:0] layer0_N85_wire = {M0[38], M0[35], M0[33], M0[18], M0[4], M0[0]};
layer0_N85 layer0_N85_inst (.M0(layer0_N85_wire), .M1(M1[85:85]));

wire [5:0] layer0_N86_wire = {M0[41], M0[36], M0[31], M0[12], M0[7], M0[6]};
layer0_N86 layer0_N86_inst (.M0(layer0_N86_wire), .M1(M1[86:86]));

wire [5:0] layer0_N87_wire = {M0[34], M0[24], M0[21], M0[18], M0[8], M0[3]};
layer0_N87 layer0_N87_inst (.M0(layer0_N87_wire), .M1(M1[87:87]));

wire [5:0] layer0_N88_wire = {M0[43], M0[29], M0[26], M0[21], M0[16], M0[7]};
layer0_N88 layer0_N88_inst (.M0(layer0_N88_wire), .M1(M1[88:88]));

wire [5:0] layer0_N89_wire = {M0[46], M0[20], M0[16], M0[9], M0[7], M0[0]};
layer0_N89 layer0_N89_inst (.M0(layer0_N89_wire), .M1(M1[89:89]));

wire [5:0] layer0_N90_wire = {M0[43], M0[31], M0[21], M0[14], M0[9], M0[5]};
layer0_N90 layer0_N90_inst (.M0(layer0_N90_wire), .M1(M1[90:90]));

wire [5:0] layer0_N91_wire = {M0[45], M0[44], M0[39], M0[22], M0[13], M0[4]};
layer0_N91 layer0_N91_inst (.M0(layer0_N91_wire), .M1(M1[91:91]));

wire [5:0] layer0_N92_wire = {M0[47], M0[38], M0[31], M0[20], M0[19], M0[6]};
layer0_N92 layer0_N92_inst (.M0(layer0_N92_wire), .M1(M1[92:92]));

wire [5:0] layer0_N93_wire = {M0[40], M0[35], M0[30], M0[27], M0[23], M0[14]};
layer0_N93 layer0_N93_inst (.M0(layer0_N93_wire), .M1(M1[93:93]));

wire [5:0] layer0_N94_wire = {M0[46], M0[39], M0[38], M0[27], M0[19], M0[1]};
layer0_N94 layer0_N94_inst (.M0(layer0_N94_wire), .M1(M1[94:94]));

wire [5:0] layer0_N95_wire = {M0[43], M0[32], M0[21], M0[14], M0[10], M0[9]};
layer0_N95 layer0_N95_inst (.M0(layer0_N95_wire), .M1(M1[95:95]));

wire [5:0] layer0_N96_wire = {M0[47], M0[42], M0[39], M0[38], M0[12], M0[5]};
layer0_N96 layer0_N96_inst (.M0(layer0_N96_wire), .M1(M1[96:96]));

wire [5:0] layer0_N97_wire = {M0[30], M0[29], M0[19], M0[13], M0[12], M0[1]};
layer0_N97 layer0_N97_inst (.M0(layer0_N97_wire), .M1(M1[97:97]));

wire [5:0] layer0_N98_wire = {M0[46], M0[39], M0[35], M0[29], M0[23], M0[16]};
layer0_N98 layer0_N98_inst (.M0(layer0_N98_wire), .M1(M1[98:98]));

wire [5:0] layer0_N99_wire = {M0[41], M0[30], M0[28], M0[25], M0[13], M0[6]};
layer0_N99 layer0_N99_inst (.M0(layer0_N99_wire), .M1(M1[99:99]));

wire [5:0] layer0_N100_wire = {M0[43], M0[42], M0[39], M0[35], M0[33], M0[12]};
layer0_N100 layer0_N100_inst (.M0(layer0_N100_wire), .M1(M1[100:100]));

wire [5:0] layer0_N101_wire = {M0[43], M0[23], M0[10], M0[8], M0[5], M0[1]};
layer0_N101 layer0_N101_inst (.M0(layer0_N101_wire), .M1(M1[101:101]));

wire [5:0] layer0_N102_wire = {M0[38], M0[36], M0[32], M0[17], M0[4], M0[3]};
layer0_N102 layer0_N102_inst (.M0(layer0_N102_wire), .M1(M1[102:102]));

wire [5:0] layer0_N103_wire = {M0[42], M0[30], M0[25], M0[21], M0[20], M0[15]};
layer0_N103 layer0_N103_inst (.M0(layer0_N103_wire), .M1(M1[103:103]));

wire [5:0] layer0_N104_wire = {M0[42], M0[41], M0[30], M0[27], M0[18], M0[8]};
layer0_N104 layer0_N104_inst (.M0(layer0_N104_wire), .M1(M1[104:104]));

wire [5:0] layer0_N105_wire = {M0[25], M0[24], M0[22], M0[18], M0[6], M0[3]};
layer0_N105 layer0_N105_inst (.M0(layer0_N105_wire), .M1(M1[105:105]));

wire [5:0] layer0_N106_wire = {M0[41], M0[36], M0[32], M0[18], M0[8], M0[0]};
layer0_N106 layer0_N106_inst (.M0(layer0_N106_wire), .M1(M1[106:106]));

wire [5:0] layer0_N107_wire = {M0[45], M0[37], M0[17], M0[6], M0[3], M0[0]};
layer0_N107 layer0_N107_inst (.M0(layer0_N107_wire), .M1(M1[107:107]));

wire [5:0] layer0_N108_wire = {M0[30], M0[19], M0[15], M0[13], M0[10], M0[4]};
layer0_N108 layer0_N108_inst (.M0(layer0_N108_wire), .M1(M1[108:108]));

wire [5:0] layer0_N109_wire = {M0[38], M0[32], M0[12], M0[11], M0[3], M0[2]};
layer0_N109 layer0_N109_inst (.M0(layer0_N109_wire), .M1(M1[109:109]));

wire [5:0] layer0_N110_wire = {M0[47], M0[43], M0[36], M0[30], M0[21], M0[6]};
layer0_N110 layer0_N110_inst (.M0(layer0_N110_wire), .M1(M1[110:110]));

wire [5:0] layer0_N111_wire = {M0[39], M0[37], M0[26], M0[18], M0[17], M0[12]};
layer0_N111 layer0_N111_inst (.M0(layer0_N111_wire), .M1(M1[111:111]));

wire [5:0] layer0_N112_wire = {M0[45], M0[36], M0[33], M0[32], M0[30], M0[9]};
layer0_N112 layer0_N112_inst (.M0(layer0_N112_wire), .M1(M1[112:112]));

wire [5:0] layer0_N113_wire = {M0[39], M0[37], M0[34], M0[29], M0[4], M0[2]};
layer0_N113 layer0_N113_inst (.M0(layer0_N113_wire), .M1(M1[113:113]));

wire [5:0] layer0_N114_wire = {M0[33], M0[30], M0[22], M0[15], M0[13], M0[9]};
layer0_N114 layer0_N114_inst (.M0(layer0_N114_wire), .M1(M1[114:114]));

wire [5:0] layer0_N115_wire = {M0[47], M0[44], M0[43], M0[24], M0[13], M0[9]};
layer0_N115 layer0_N115_inst (.M0(layer0_N115_wire), .M1(M1[115:115]));

wire [5:0] layer0_N116_wire = {M0[45], M0[31], M0[23], M0[15], M0[8], M0[5]};
layer0_N116 layer0_N116_inst (.M0(layer0_N116_wire), .M1(M1[116:116]));

wire [5:0] layer0_N117_wire = {M0[35], M0[32], M0[28], M0[19], M0[13], M0[11]};
layer0_N117 layer0_N117_inst (.M0(layer0_N117_wire), .M1(M1[117:117]));

wire [5:0] layer0_N118_wire = {M0[41], M0[39], M0[37], M0[34], M0[24], M0[6]};
layer0_N118 layer0_N118_inst (.M0(layer0_N118_wire), .M1(M1[118:118]));

wire [5:0] layer0_N119_wire = {M0[35], M0[33], M0[31], M0[18], M0[13], M0[0]};
layer0_N119 layer0_N119_inst (.M0(layer0_N119_wire), .M1(M1[119:119]));

wire [5:0] layer0_N120_wire = {M0[29], M0[28], M0[20], M0[16], M0[15], M0[14]};
layer0_N120 layer0_N120_inst (.M0(layer0_N120_wire), .M1(M1[120:120]));

wire [5:0] layer0_N121_wire = {M0[45], M0[41], M0[35], M0[32], M0[11], M0[4]};
layer0_N121 layer0_N121_inst (.M0(layer0_N121_wire), .M1(M1[121:121]));

wire [5:0] layer0_N122_wire = {M0[45], M0[40], M0[38], M0[34], M0[14], M0[5]};
layer0_N122 layer0_N122_inst (.M0(layer0_N122_wire), .M1(M1[122:122]));

wire [5:0] layer0_N123_wire = {M0[46], M0[38], M0[33], M0[22], M0[11], M0[5]};
layer0_N123 layer0_N123_inst (.M0(layer0_N123_wire), .M1(M1[123:123]));

wire [5:0] layer0_N124_wire = {M0[44], M0[25], M0[24], M0[23], M0[16], M0[15]};
layer0_N124 layer0_N124_inst (.M0(layer0_N124_wire), .M1(M1[124:124]));

wire [5:0] layer0_N125_wire = {M0[44], M0[37], M0[34], M0[26], M0[21], M0[20]};
layer0_N125 layer0_N125_inst (.M0(layer0_N125_wire), .M1(M1[125:125]));

wire [5:0] layer0_N126_wire = {M0[45], M0[43], M0[30], M0[22], M0[17], M0[5]};
layer0_N126 layer0_N126_inst (.M0(layer0_N126_wire), .M1(M1[126:126]));

wire [5:0] layer0_N127_wire = {M0[45], M0[44], M0[41], M0[15], M0[7], M0[4]};
layer0_N127 layer0_N127_inst (.M0(layer0_N127_wire), .M1(M1[127:127]));

wire [5:0] layer0_N128_wire = {M0[44], M0[43], M0[30], M0[6], M0[3], M0[1]};
layer0_N128 layer0_N128_inst (.M0(layer0_N128_wire), .M1(M1[128:128]));

wire [5:0] layer0_N129_wire = {M0[45], M0[35], M0[27], M0[14], M0[10], M0[7]};
layer0_N129 layer0_N129_inst (.M0(layer0_N129_wire), .M1(M1[129:129]));

wire [5:0] layer0_N130_wire = {M0[45], M0[17], M0[14], M0[12], M0[11], M0[2]};
layer0_N130 layer0_N130_inst (.M0(layer0_N130_wire), .M1(M1[130:130]));

wire [5:0] layer0_N131_wire = {M0[38], M0[25], M0[22], M0[21], M0[18], M0[11]};
layer0_N131 layer0_N131_inst (.M0(layer0_N131_wire), .M1(M1[131:131]));

wire [5:0] layer0_N132_wire = {M0[46], M0[30], M0[29], M0[20], M0[4], M0[2]};
layer0_N132 layer0_N132_inst (.M0(layer0_N132_wire), .M1(M1[132:132]));

wire [5:0] layer0_N133_wire = {M0[40], M0[31], M0[30], M0[21], M0[11], M0[0]};
layer0_N133 layer0_N133_inst (.M0(layer0_N133_wire), .M1(M1[133:133]));

wire [5:0] layer0_N134_wire = {M0[42], M0[27], M0[20], M0[18], M0[16], M0[6]};
layer0_N134 layer0_N134_inst (.M0(layer0_N134_wire), .M1(M1[134:134]));

wire [5:0] layer0_N135_wire = {M0[42], M0[37], M0[23], M0[15], M0[14], M0[2]};
layer0_N135 layer0_N135_inst (.M0(layer0_N135_wire), .M1(M1[135:135]));

wire [5:0] layer0_N136_wire = {M0[37], M0[36], M0[16], M0[8], M0[1], M0[0]};
layer0_N136 layer0_N136_inst (.M0(layer0_N136_wire), .M1(M1[136:136]));

wire [5:0] layer0_N137_wire = {M0[45], M0[28], M0[21], M0[14], M0[13], M0[1]};
layer0_N137 layer0_N137_inst (.M0(layer0_N137_wire), .M1(M1[137:137]));

wire [5:0] layer0_N138_wire = {M0[46], M0[30], M0[19], M0[18], M0[17], M0[6]};
layer0_N138 layer0_N138_inst (.M0(layer0_N138_wire), .M1(M1[138:138]));

wire [5:0] layer0_N139_wire = {M0[40], M0[37], M0[31], M0[15], M0[12], M0[1]};
layer0_N139 layer0_N139_inst (.M0(layer0_N139_wire), .M1(M1[139:139]));

wire [5:0] layer0_N140_wire = {M0[46], M0[45], M0[21], M0[8], M0[4], M0[0]};
layer0_N140 layer0_N140_inst (.M0(layer0_N140_wire), .M1(M1[140:140]));

wire [5:0] layer0_N141_wire = {M0[39], M0[36], M0[25], M0[11], M0[4], M0[3]};
layer0_N141 layer0_N141_inst (.M0(layer0_N141_wire), .M1(M1[141:141]));

wire [5:0] layer0_N142_wire = {M0[47], M0[42], M0[35], M0[24], M0[3], M0[0]};
layer0_N142 layer0_N142_inst (.M0(layer0_N142_wire), .M1(M1[142:142]));

wire [5:0] layer0_N143_wire = {M0[37], M0[25], M0[19], M0[14], M0[10], M0[1]};
layer0_N143 layer0_N143_inst (.M0(layer0_N143_wire), .M1(M1[143:143]));

wire [5:0] layer0_N144_wire = {M0[41], M0[25], M0[24], M0[15], M0[14], M0[3]};
layer0_N144 layer0_N144_inst (.M0(layer0_N144_wire), .M1(M1[144:144]));

endmodule